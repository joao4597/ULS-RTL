// Simple Dual-Port Block RAM with One Clock
// File: simple_dual_one_clock.v

/**
 * GENERAL DESCRIPTION:
 *
 * -16 bit by 512 lines RAM that holds the 512 coefficients of a Band Pass filter
 * -FPass_1 -> 15KHz || FCut_1 -> 18KHz || FCut_2 -> 32KHz || FPass_2 -> 35 KHz
 *
 *
 * CONSTRAINTS:
 *
 *
 */


module rx_BRAM_16_512_band_pass (clk, rrx_rst, ena,enb,wea,addra,addrb,dia,dob);

  input                clk    ;  //clock
  input                rrx_rst;
  input                ena    ;  //enable
  input                enb    ;  //enable read
  input                wea    ;  //write enable
  input          [8:0] addra  ;  //write address
  input          [8:0] addrb  ;  //read addr
  input  signed [15:0] dia    ;  //data in
  output signed [15:0] dob    ;  //data out

  reg signed [15:0] ram [511:0];
  reg signed [15:0] doa         ;
  reg signed [15:0] dob         ;

  integer i;

  //set iniial value of memories to zero
  initial begin
    ram[0] = 0;
    ram[1] = 1;
    ram[2] = 0;
    ram[3] = 0;
    ram[4] = 0;
    ram[5] = 0;
    ram[6] = 0;
    ram[7] = 0;
    ram[8] = 0;
    ram[9] = 0;
    ram[10] = 0;
    ram[11] = 0;
    ram[12] = 0;
    ram[13] = 0;
    ram[14] = 0;
    ram[15] = 0;
    ram[16] = 0;
    ram[17] = 0;
    ram[18] = 0;
    ram[19] = 0;
    ram[20] = 0;
    ram[21] = 0;
    ram[22] = 0;
    ram[23] = 0;
    ram[24] = 0;
    ram[25] = 0;
    ram[26] = 0;
    ram[27] = 0;
    ram[28] = 0;
    ram[29] = 0;
    ram[30] = 0;
    ram[31] = 0;
    ram[32] = 0;
    ram[33] = 0;
    ram[34] = 0;
    ram[35] = 0;
    ram[36] = 0;
    ram[37] = 0;
    ram[38] = 0;
    ram[39] = 0;
    ram[40] = 0;
    ram[41] = 0;
    ram[42] = 0;
    ram[43] = 0;
    ram[44] = 0;
    ram[45] = 0;
    ram[46] = 0;
    ram[47] = 0;
    ram[48] = 0;
    ram[49] = 0;
    ram[50] = 0;
    ram[51] = 1;
    ram[52] = 0;
    ram[53] = 0;
    ram[54] = 0;
    ram[55] = -1;
    ram[56] = -1;
    ram[57] = 0;
    ram[58] = 0;
    ram[59] = 0;
    ram[60] = 0;
    ram[61] = 0;
    ram[62] = 0;
    ram[63] = 0;
    ram[64] = 1;
    ram[65] = 1;
    ram[66] = 1;
    ram[67] = 0;
    ram[68] = 0;
    ram[69] = -1;
    ram[70] = -1;
    ram[71] = -1;
    ram[72] = 0;
    ram[73] = 0;
    ram[74] = 0;
    ram[75] = 0;
    ram[76] = 0;
    ram[77] = 0;
    ram[78] = 0;
    ram[79] = 1;
    ram[80] = 1;
    ram[81] = 1;
    ram[82] = 0;
    ram[83] = -1;
    ram[84] = -1;
    ram[85] = -1;
    ram[86] = 0;
    ram[87] = 0;
    ram[88] = 0;
    ram[89] = 0;
    ram[90] = -1;
    ram[91] = -1;
    ram[92] = 0;
    ram[93] = 1;
    ram[94] = 2;
    ram[95] = 2;
    ram[96] = 1;
    ram[97] = 0;
    ram[98] = -1;
    ram[99] = -1;
    ram[100] = -1;
    ram[101] = 0;
    ram[102] = 0;
    ram[103] = 0;
    ram[104] = -1;
    ram[105] = -1;
    ram[106] = -1;
    ram[107] = 1;
    ram[108] = 2;
    ram[109] = 2;
    ram[110] = 2;
    ram[111] = 1;
    ram[112] = -1;
    ram[113] = -1;
    ram[114] = -1;
    ram[115] = 0;
    ram[116] = 0;
    ram[117] = 0;
    ram[118] = -1;
    ram[119] = -2;
    ram[120] = -1;
    ram[121] = 0;
    ram[122] = 1;
    ram[123] = 3;
    ram[124] = 3;
    ram[125] = 2;
    ram[126] = 0;
    ram[127] = -1;
    ram[128] = -1;
    ram[129] = -1;
    ram[130] = 0;
    ram[131] = 0;
    ram[132] = -1;
    ram[133] = -2;
    ram[134] = -2;
    ram[135] = -2;
    ram[136] = 0;
    ram[137] = 2;
    ram[138] = 3;
    ram[139] = 3;
    ram[140] = 1;
    ram[141] = 0;
    ram[142] = -1;
    ram[143] = -1;
    ram[144] = 0;
    ram[145] = 0;
    ram[146] = 0;
    ram[147] = -2;
    ram[148] = -3;
    ram[149] = -3;
    ram[150] = -1;
    ram[151] = 1;
    ram[152] = 4;
    ram[153] = 4;
    ram[154] = 3;
    ram[155] = 1;
    ram[156] = -1;
    ram[157] = -1;
    ram[158] = 0;
    ram[159] = 1;
    ram[160] = 0;
    ram[161] = -1;
    ram[162] = -4;
    ram[163] = -5;
    ram[164] = -4;
    ram[165] = -1;
    ram[166] = 3;
    ram[167] = 5;
    ram[168] = 4;
    ram[169] = 2;
    ram[170] = 0;
    ram[171] = -1;
    ram[172] = 0;
    ram[173] = 2;
    ram[174] = 2;
    ram[175] = 0;
    ram[176] = -3;
    ram[177] = -6;
    ram[178] = -6;
    ram[179] = -4;
    ram[180] = 1;
    ram[181] = 4;
    ram[182] = 6;
    ram[183] = 4;
    ram[184] = 1;
    ram[185] = 0;
    ram[186] = 0;
    ram[187] = 2;
    ram[188] = 3;
    ram[189] = 2;
    ram[190] = -2;
    ram[191] = -6;
    ram[192] = -9;
    ram[193] = -7;
    ram[194] = -3;
    ram[195] = 3;
    ram[196] = 6;
    ram[197] = 6;
    ram[198] = 3;
    ram[199] = 0;
    ram[200] = 0;
    ram[201] = 3;
    ram[202] = 5;
    ram[203] = 5;
    ram[204] = 1;
    ram[205] = -5;
    ram[206] = -11;
    ram[207] = -12;
    ram[208] = -8;
    ram[209] = -1;
    ram[210] = 5;
    ram[211] = 7;
    ram[212] = 5;
    ram[213] = 1;
    ram[214] = 0;
    ram[215] = 3;
    ram[216] = 8;
    ram[217] = 10;
    ram[218] = 7;
    ram[219] = -1;
    ram[220] = -12;
    ram[221] = -18;
    ram[222] = -16;
    ram[223] = -8;
    ram[224] = 2;
    ram[225] = 8;
    ram[226] = 8;
    ram[227] = 3;
    ram[228] = -1;
    ram[229] = 2;
    ram[230] = 10;
    ram[231] = 18;
    ram[232] = 19;
    ram[233] = 9;
    ram[234] = -9;
    ram[235] = -25;
    ram[236] = -31;
    ram[237] = -23;
    ram[238] = -7;
    ram[239] = 8;
    ram[240] = 12;
    ram[241] = 5;
    ram[242] = -4;
    ram[243] = -3;
    ram[244] = 13;
    ram[245] = 39;
    ram[246] = 57;
    ram[247] = 49;
    ram[248] = 10;
    ram[249] = -50;
    ram[250] = -103;
    ram[251] = -119;
    ram[252] = -83;
    ram[253] = -5;
    ram[254] = 82;
    ram[255] = 139;
    ram[256] = 139;
    ram[257] = 82;
    ram[258] = -5;
    ram[259] = -83;
    ram[260] = -119;
    ram[261] = -103;
    ram[262] = -50;
    ram[263] = 10;
    ram[264] = 49;
    ram[265] = 57;
    ram[266] = 39;
    ram[267] = 13;
    ram[268] = -3;
    ram[269] = -4;
    ram[270] = 5;
    ram[271] = 12;
    ram[272] = 8;
    ram[273] = -7;
    ram[274] = -23;
    ram[275] = -31;
    ram[276] = -25;
    ram[277] = -9;
    ram[278] = 9;
    ram[279] = 19;
    ram[280] = 18;
    ram[281] = 10;
    ram[282] = 2;
    ram[283] = -1;
    ram[284] = 3;
    ram[285] = 8;
    ram[286] = 8;
    ram[287] = 2;
    ram[288] = -8;
    ram[289] = -16;
    ram[290] = -18;
    ram[291] = -12;
    ram[292] = -1;
    ram[293] = 7;
    ram[294] = 10;
    ram[295] = 8;
    ram[296] = 3;
    ram[297] = 0;
    ram[298] = 1;
    ram[299] = 5;
    ram[300] = 7;
    ram[301] = 5;
    ram[302] = -1;
    ram[303] = -8;
    ram[304] = -12;
    ram[305] = -11;
    ram[306] = -5;
    ram[307] = 1;
    ram[308] = 5;
    ram[309] = 5;
    ram[310] = 3;
    ram[311] = 0;
    ram[312] = 0;
    ram[313] = 3;
    ram[314] = 6;
    ram[315] = 6;
    ram[316] = 3;
    ram[317] = -3;
    ram[318] = -7;
    ram[319] = -9;
    ram[320] = -6;
    ram[321] = -2;
    ram[322] = 2;
    ram[323] = 3;
    ram[324] = 2;
    ram[325] = 0;
    ram[326] = 0;
    ram[327] = 1;
    ram[328] = 4;
    ram[329] = 6;
    ram[330] = 4;
    ram[331] = 1;
    ram[332] = -4;
    ram[333] = -6;
    ram[334] = -6;
    ram[335] = -3;
    ram[336] = 0;
    ram[337] = 2;
    ram[338] = 2;
    ram[339] = 0;
    ram[340] = -1;
    ram[341] = 0;
    ram[342] = 2;
    ram[343] = 4;
    ram[344] = 5;
    ram[345] = 3;
    ram[346] = -1;
    ram[347] = -4;
    ram[348] = -5;
    ram[349] = -4;
    ram[350] = -1;
    ram[351] = 0;
    ram[352] = 1;
    ram[353] = 0;
    ram[354] = -1;
    ram[355] = -1;
    ram[356] = 1;
    ram[357] = 3;
    ram[358] = 4;
    ram[359] = 4;
    ram[360] = 1;
    ram[361] = -1;
    ram[362] = -3;
    ram[363] = -3;
    ram[364] = -2;
    ram[365] = 0;
    ram[366] = 0;
    ram[367] = 0;
    ram[368] = -1;
    ram[369] = -1;
    ram[370] = 0;
    ram[371] = 1;
    ram[372] = 3;
    ram[373] = 3;
    ram[374] = 2;
    ram[375] = 0;
    ram[376] = -2;
    ram[377] = -2;
    ram[378] = -2;
    ram[379] = -1;
    ram[380] = 0;
    ram[381] = 0;
    ram[382] = -1;
    ram[383] = -1;
    ram[384] = -1;
    ram[385] = 0;
    ram[386] = 2;
    ram[387] = 3;
    ram[388] = 3;
    ram[389] = 1;
    ram[390] = 0;
    ram[391] = -1;
    ram[392] = -2;
    ram[393] = -1;
    ram[394] = 0;
    ram[395] = 0;
    ram[396] = 0;
    ram[397] = -1;
    ram[398] = -1;
    ram[399] = -1;
    ram[400] = 1;
    ram[401] = 2;
    ram[402] = 2;
    ram[403] = 2;
    ram[404] = 1;
    ram[405] = -1;
    ram[406] = -1;
    ram[407] = -1;
    ram[408] = 0;
    ram[409] = 0;
    ram[410] = 0;
    ram[411] = -1;
    ram[412] = -1;
    ram[413] = -1;
    ram[414] = 0;
    ram[415] = 1;
    ram[416] = 2;
    ram[417] = 2;
    ram[418] = 1;
    ram[419] = 0;
    ram[420] = -1;
    ram[421] = -1;
    ram[422] = 0;
    ram[423] = 0;
    ram[424] = 0;
    ram[425] = 0;
    ram[426] = -1;
    ram[427] = -1;
    ram[428] = -1;
    ram[429] = 0;
    ram[430] = 1;
    ram[431] = 1;
    ram[432] = 1;
    ram[433] = 0;
    ram[434] = 0;
    ram[435] = 0;
    ram[436] = 0;
    ram[437] = 0;
    ram[438] = 0;
    ram[439] = 0;
    ram[440] = -1;
    ram[441] = -1;
    ram[442] = -1;
    ram[443] = 0;
    ram[444] = 0;
    ram[445] = 1;
    ram[446] = 1;
    ram[447] = 1;
    ram[448] = 0;
    ram[449] = 0;
    ram[450] = 0;
    ram[451] = 0;
    ram[452] = 0;
    ram[453] = 0;
    ram[454] = 0;
    ram[455] = -1;
    ram[456] = -1;
    ram[457] = 0;
    ram[458] = 0;
    ram[459] = 0;
    ram[460] = 1;
    ram[461] = 0;
    ram[462] = 0;
    ram[463] = 0;
    ram[464] = 0;
    ram[465] = 0;
    ram[466] = 0;
    ram[467] = 0;
    ram[468] = 0;
    ram[469] = 0;
    ram[470] = 0;
    ram[471] = 0;
    ram[472] = 0;
    ram[473] = 0;
    ram[474] = 0;
    ram[475] = 0;
    ram[476] = 0;
    ram[477] = 0;
    ram[478] = 0;
    ram[479] = 0;
    ram[480] = 0;
    ram[481] = 0;
    ram[482] = 0;
    ram[483] = 0;
    ram[484] = 0;
    ram[485] = 0;
    ram[486] = 0;
    ram[487] = 0;
    ram[488] = 0;
    ram[489] = 0;
    ram[490] = 0;
    ram[491] = 0;
    ram[492] = 0;
    ram[493] = 0;
    ram[494] = 0;
    ram[495] = 0;
    ram[496] = 0;
    ram[497] = 0;
    ram[498] = 0;
    ram[499] = 0;
    ram[500] = 0;
    ram[501] = 0;
    ram[502] = 0;
    ram[503] = 0;
    ram[504] = 0;
    ram[505] = 0;
    ram[506] = 0;
    ram[507] = 0;
    ram[508] = 0;
    ram[509] = 0;
    ram[510] = 1;
    ram[511] = 0;

    dob = ram[511];
  end

  always @(posedge clk) begin
   if (ena) begin
      if (wea)
          ram[addra] <= dia;
   end
  end

  always @(posedge clk) begin
    if (rrx_rst) begin
      dob <= ram[511];
    end else begin
      if (enb) begin
        dob <= ram[addrb];
      end
    end
  end

endmodule
