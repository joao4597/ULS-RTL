// Simple Dual-Port Block RAM with One Clock
// File: simple_dual_one_clock.v


//16 by 256
module rx_BRAM_16_256_binary_sequences (clk,ena,enb,wea,addra,addrb,dia,dob);
  
  input         clk  ;  //clock
  input         ena  ;  //enable
  input         enb  ;  //enable read
  input         wea  ;  //write enable
  input  [7:0]  addra;  //write address
  input  [7:0]  addrb;  //read addr
  input  [15:0] dia  ;  //data in
  output [15:0] dob  ;  //data out
  
  reg [15:0] ram [255:0];
  reg [15:0] doa        ;
  reg [15:0] dob        ;
  
  //Initalize the ram with the 16 possible binary sequences
  //each collum represents a sequence
  initial begin
    ram[0]   = 16'b0110001001101011;
    ram[1]   = 16'b1000111011001010;
    ram[2]   = 16'b1000011101100101;
    ram[3]   = 16'b0011110001001101;
    ram[4]   = 16'b0101111000100110;
    ram[5]   = 16'b0010111100010011;
    ram[6]   = 16'b1010100001110110;
    ram[7]   = 16'b1001010000111011;
    ram[8]   = 16'b1100101000011101;
    ram[9]   = 16'b1110010100001110;
    ram[10]  = 16'b0100110101111000;
    ram[11]  = 16'b1101100101000011;
    ram[12]  = 16'b0001001101011110;
    ram[13]  = 16'b0000100110101111;
    ram[14]  = 16'b0100010011010111;
    ram[15]  = 16'b0110001001101011;
    ram[16]  = 16'b1000111011001010;
    ram[17]  = 16'b1000011101100101;
    ram[18]  = 16'b1100001110110010;
    ram[19]  = 16'b1010000111011001;
    ram[20]  = 16'b1101000011101100;
    ram[21]  = 16'b1010100001110110;
    ram[22]  = 16'b1001010000111011;
    ram[23]  = 16'b1100101000011101;
    ram[24]  = 16'b0001101011110001;
    ram[25]  = 16'b0100110101111000;
    ram[26]  = 16'b1101100101000011;
    ram[27]  = 16'b0001001101011110;
    ram[28]  = 16'b0000100110101111;
    ram[29]  = 16'b0100010011010111;
    ram[30]  = 16'b0110001001101011;
    ram[31]  = 16'b1000111011001010;
    ram[32]  = 16'b0111100010011010;
    ram[33]  = 16'b1100001110110010;
    ram[34]  = 16'b0101111000100110;
    ram[35]  = 16'b0010111100010011;
    ram[36]  = 16'b1010100001110110;
    ram[37]  = 16'b1001010000111011;
    ram[38]  = 16'b1100101000011101;
    ram[39]  = 16'b1110010100001110;
    ram[40]  = 16'b1011001010000111;
    ram[41]  = 16'b0010011010111100;
    ram[42]  = 16'b1110110010100001;
    ram[43]  = 16'b0000100110101111;
    ram[44]  = 16'b1011101100101000;
    ram[45]  = 16'b0110001001101011;
    ram[46]  = 16'b1000111011001010;
    ram[47]  = 16'b0111100010011010;
    ram[48]  = 16'b1100001110110010;
    ram[49]  = 16'b1010000111011001;
    ram[50]  = 16'b1101000011101100;
    ram[51]  = 16'b0101011110001001;
    ram[52]  = 16'b0110101111000100;
    ram[53]  = 16'b0011010111100010;
    ram[54]  = 16'b0001101011110001;
    ram[55]  = 16'b0100110101111000;
    ram[56]  = 16'b1101100101000011;
    ram[57]  = 16'b1110110010100001;
    ram[58]  = 16'b0000100110101111;
    ram[59]  = 16'b0100010011010111;
    ram[60]  = 16'b0110001001101011;
    ram[61]  = 16'b1000111011001010;
    ram[62]  = 16'b0111100010011010;
    ram[63]  = 16'b1100001110110010;
    ram[64]  = 16'b0101111000100110;
    ram[65]  = 16'b1101000011101100;
    ram[66]  = 16'b1010100001110110;
    ram[67]  = 16'b0110101111000100;
    ram[68]  = 16'b0011010111100010;
    ram[69]  = 16'b1110010100001110;
    ram[70]  = 16'b1011001010000111;
    ram[71]  = 16'b0010011010111100;
    ram[72]  = 16'b0001001101011110;
    ram[73]  = 16'b1111011001010000;
    ram[74]  = 16'b0100010011010111;
    ram[75]  = 16'b1001110110010100;
    ram[76]  = 16'b1000111011001010;
    ram[77]  = 16'b1000011101100101;
    ram[78]  = 16'b1100001110110010;
    ram[79]  = 16'b1010000111011001;
    ram[80]  = 16'b1101000011101100;
    ram[81]  = 16'b0101011110001001;
    ram[82]  = 16'b1001010000111011;
    ram[83]  = 16'b1100101000011101;
    ram[84]  = 16'b1110010100001110;
    ram[85]  = 16'b1011001010000111;
    ram[86]  = 16'b0010011010111100;
    ram[87]  = 16'b0001001101011110;
    ram[88]  = 16'b1111011001010000;
    ram[89]  = 16'b1011101100101000;
    ram[90]  = 16'b0110001001101011;
    ram[91]  = 16'b1000111011001010;
    ram[92]  = 16'b1000011101100101;
    ram[93]  = 16'b1100001110110010;
    ram[94]  = 16'b0101111000100110;
    ram[95]  = 16'b1101000011101100;
    ram[96]  = 16'b1010100001110110;
    ram[97]  = 16'b1001010000111011;
    ram[98]  = 16'b0011010111100010;
    ram[99]  = 16'b0001101011110001;
    ram[100] = 16'b1011001010000111;
    ram[101] = 16'b0010011010111100;
    ram[102] = 16'b1110110010100001;
    ram[103] = 16'b0000100110101111;
    ram[104] = 16'b1011101100101000;
    ram[105] = 16'b0110001001101011;
    ram[106] = 16'b0111000100110101;
    ram[107] = 16'b1000011101100101;
    ram[108] = 16'b0011110001001101;
    ram[109] = 16'b1010000111011001;
    ram[110] = 16'b0010111100010011;
    ram[111] = 16'b0101011110001001;
    ram[112] = 16'b0110101111000100;
    ram[113] = 16'b1100101000011101;
    ram[114] = 16'b0001101011110001;
    ram[115] = 16'b0100110101111000;
    ram[116] = 16'b1101100101000011;
    ram[117] = 16'b0001001101011110;
    ram[118] = 16'b1111011001010000;
    ram[119] = 16'b1011101100101000;
    ram[120] = 16'b0110001001101011;
    ram[121] = 16'b1000111011001010;
    ram[122] = 16'b0111100010011010;
    ram[123] = 16'b0011110001001101;
    ram[124] = 16'b0101111000100110;
    ram[125] = 16'b1101000011101100;
    ram[126] = 16'b1010100001110110;
    ram[127] = 16'b0110101111000100;
    ram[128] = 16'b0011010111100010;
    ram[129] = 16'b1110010100001110;
    ram[130] = 16'b1011001010000111;
    ram[131] = 16'b1101100101000011;
    ram[132] = 16'b0001001101011110;
    ram[133] = 16'b0000100110101111;
    ram[134] = 16'b1011101100101000;
    ram[135] = 16'b1001110110010100;
    ram[136] = 16'b1000111011001010;
    ram[137] = 16'b1000011101100101;
    ram[138] = 16'b0011110001001101;
    ram[139] = 16'b0101111000100110;
    ram[140] = 16'b0010111100010011;
    ram[141] = 16'b1010100001110110;
    ram[142] = 16'b1001010000111011;
    ram[143] = 16'b0011010111100010;
    ram[144] = 16'b1110010100001110;
    ram[145] = 16'b1011001010000111;
    ram[146] = 16'b0010011010111100;
    ram[147] = 16'b0001001101011110;
    ram[148] = 16'b0000100110101111;
    ram[149] = 16'b0100010011010111;
    ram[150] = 16'b1001110110010100;
    ram[151] = 16'b0111000100110101;
    ram[152] = 16'b0111100010011010;
    ram[153] = 16'b0011110001001101;
    ram[154] = 16'b1010000111011001;
    ram[155] = 16'b0010111100010011;
    ram[156] = 16'b1010100001110110;
    ram[157] = 16'b1001010000111011;
    ram[158] = 16'b1100101000011101;
    ram[159] = 16'b0001101011110001;
    ram[160] = 16'b1011001010000111;
    ram[161] = 16'b0010011010111100;
    ram[162] = 16'b1110110010100001;
    ram[163] = 16'b1111011001010000;
    ram[164] = 16'b1011101100101000;
    ram[165] = 16'b1001110110010100;
    ram[166] = 16'b0111000100110101;
    ram[167] = 16'b1000011101100101;
    ram[168] = 16'b1100001110110010;
    ram[169] = 16'b0101111000100110;
    ram[170] = 16'b1101000011101100;
    ram[171] = 16'b1010100001110110;
    ram[172] = 16'b1001010000111011;
    ram[173] = 16'b1100101000011101;
    ram[174] = 16'b1110010100001110;
    ram[175] = 16'b0100110101111000;
    ram[176] = 16'b0010011010111100;
    ram[177] = 16'b0001001101011110;
    ram[178] = 16'b0000100110101111;
    ram[179] = 16'b1011101100101000;
    ram[180] = 16'b1001110110010100;
    ram[181] = 16'b0111000100110101;
    ram[182] = 16'b1000011101100101;
    ram[183] = 16'b0011110001001101;
    ram[184] = 16'b0101111000100110;
    ram[185] = 16'b1101000011101100;
    ram[186] = 16'b1010100001110110;
    ram[187] = 16'b0110101111000100;
    ram[188] = 16'b1100101000011101;
    ram[189] = 16'b0001101011110001;
    ram[190] = 16'b1011001010000111;
    ram[191] = 16'b1101100101000011;
    ram[192] = 16'b0001001101011110;
    ram[193] = 16'b1111011001010000;
    ram[194] = 16'b1011101100101000;
    ram[195] = 16'b0110001001101011;
    ram[196] = 16'b1000111011001010;
    ram[197] = 16'b0111100010011010;
    ram[198] = 16'b1100001110110010;
    ram[199] = 16'b0101111000100110;
    ram[200] = 16'b0010111100010011;
    ram[201] = 16'b0101011110001001;
    ram[202] = 16'b0110101111000100;
    ram[203] = 16'b0011010111100010;
    ram[204] = 16'b1110010100001110;
    ram[205] = 16'b0100110101111000;
    ram[206] = 16'b0010011010111100;
    ram[207] = 16'b1110110010100001;
    ram[208] = 16'b1111011001010000;
    ram[209] = 16'b1011101100101000;
    ram[210] = 16'b0110001001101011;
    ram[211] = 16'b1000111011001010;
    ram[212] = 16'b1000011101100101;
    ram[213] = 16'b0011110001001101;
    ram[214] = 16'b0101111000100110;
    ram[215] = 16'b1101000011101100;
    ram[216] = 16'b0101011110001001;
    ram[217] = 16'b0110101111000100;
    ram[218] = 16'b1100101000011101;
    ram[219] = 16'b0001101011110001;
    ram[220] = 16'b0100110101111000;
    ram[221] = 16'b1101100101000011;
    ram[222] = 16'b1110110010100001;
    ram[223] = 16'b0000100110101111;
    ram[224] = 16'b0100010011010111;
    ram[225] = 16'b0110001001101011;
    ram[226] = 16'b0111000100110101;
    ram[227] = 16'b0111100010011010;
    ram[228] = 16'b0011110001001101;
    ram[229] = 16'b1010000111011001;
    ram[230] = 16'b1101000011101100;
    ram[231] = 16'b1010100001110110;
    ram[232] = 16'b0110101111000100;
    ram[233] = 16'b1100101000011101;
    ram[234] = 16'b0001101011110001;
    ram[235] = 16'b0100110101111000;
    ram[236] = 16'b1101100101000011;
    ram[237] = 16'b0001001101011110;
    ram[238] = 16'b0000100110101111;
    ram[239] = 16'b0100010011010111;
    ram[240] = 16'b1001110110010100;
    ram[241] = 16'b1000111011001010;
    ram[242] = 16'b1000011101100101;
    ram[243] = 16'b0011110001001101;
    ram[244] = 16'b0101111000100110;
    ram[245] = 16'b0010111100010011;
    ram[246] = 16'b1010100001110110;
    ram[247] = 16'b0110101111000100;
    ram[248] = 16'b0011010111100010;
    ram[249] = 16'b0001101011110001;
    ram[250] = 16'b0100110101111000;
    ram[251] = 16'b0010011010111100;
    ram[252] = 16'b0001001101011110;
    ram[253] = 16'b0000100110101111;
    ram[254] = 16'b1011101100101000;
  end
  
  always @(posedge clk) begin 
   if (ena) begin
      if (wea)
          ram[addra] <= dia;
   end
  end
    
  always @(posedge clk) begin 
    if (enb)
      dob <= ram[addrb];
  end
  
endmodule

//MODULE OBTAINED ON THE XILINX WEBSITE