// Simple Dual-Port Block RAM with One Clock
// File: simple_dual_one_clock.v


//16 by 256
module rx_BRAM_16_256 (clk,ena,enb,wea,addra,addrb,dia,dob);
  
  input         clk  ;  //clock
  input         ena  ;  //enable
  input         enb  ;  //enable read
  input         wea  ;  //write enable
  input  [7:0]  addra;  //write address
  input  [7:0]  addrb;  //read addr
  input  [15:0] dia  ;  //data in
  output [15:0] dob  ;  //data out
  
  reg [15:0] ram [255:0];
  reg [15:0] doa         ;
  reg [15:0] dob         ;
  
  //Initalize the ram with the 16 possible binary sequences
  //each collum represents a sequence
  initial begin
    ram[0]   = 0110001001101011;
    ram[1]   = 1000111011001010;
    ram[2]   = 1000011101100101;
    ram[3]   = 0011110001001101;
    ram[4]   = 0101111000100110;
    ram[5]   = 0010111100010011;
    ram[6]   = 1010100001110110;
    ram[7]   = 1001010000111011;
    ram[8]   = 1100101000011101;
    ram[9]   = 1110010100001110;
    ram[10]  = 0100110101111000;
    ram[11]  = 1101100101000011;
    ram[12]  = 0001001101011110;
    ram[13]  = 0000100110101111;
    ram[14]  = 0100010011010111;
    ram[15]  = 0110001001101011;
    ram[16]  = 1000111011001010;
    ram[17]  = 1000011101100101;
    ram[18]  = 1100001110110010;
    ram[19]  = 1010000111011001;
    ram[20]  = 1101000011101100;
    ram[21]  = 1010100001110110;
    ram[22]  = 1001010000111011;
    ram[23]  = 1100101000011101;
    ram[24]  = 0001101011110001;
    ram[25]  = 0100110101111000;
    ram[26]  = 1101100101000011;
    ram[27]  = 0001001101011110;
    ram[28]  = 0000100110101111;
    ram[29]  = 0100010011010111;
    ram[30]  = 0110001001101011;
    ram[31]  = 1000111011001010;
    ram[32]  = 0111100010011010;
    ram[33]  = 1100001110110010;
    ram[34]  = 0101111000100110;
    ram[35]  = 0010111100010011;
    ram[36]  = 1010100001110110;
    ram[37]  = 1001010000111011;
    ram[38]  = 1100101000011101;
    ram[39]  = 1110010100001110;
    ram[40]  = 1011001010000111;
    ram[41]  = 0010011010111100;
    ram[42]  = 1110110010100001;
    ram[43]  = 0000100110101111;
    ram[44]  = 1011101100101000;
    ram[45]  = 0110001001101011;
    ram[46]  = 1000111011001010;
    ram[47]  = 0111100010011010;
    ram[48]  = 1100001110110010;
    ram[49]  = 1010000111011001;
    ram[50]  = 1101000011101100;
    ram[51]  = 0101011110001001;
    ram[52]  = 0110101111000100;
    ram[53]  = 0011010111100010;
    ram[54]  = 0001101011110001;
    ram[55]  = 0100110101111000;
    ram[56]  = 1101100101000011;
    ram[57]  = 1110110010100001;
    ram[58]  = 0000100110101111;
    ram[59]  = 0100010011010111;
    ram[60]  = 0110001001101011;
    ram[61]  = 1000111011001010;
    ram[62]  = 0111100010011010;
    ram[63]  = 1100001110110010;
    ram[64]  = 0101111000100110;
    ram[65]  = 1101000011101100;
    ram[66]  = 1010100001110110;
    ram[67]  = 0110101111000100;
    ram[68]  = 0011010111100010;
    ram[69]  = 1110010100001110;
    ram[70]  = 1011001010000111;
    ram[71]  = 0010011010111100;
    ram[72]  = 0001001101011110;
    ram[73]  = 1111011001010000;
    ram[74]  = 0100010011010111;
    ram[75]  = 1001110110010100;
    ram[76]  = 1000111011001010;
    ram[77]  = 1000011101100101;
    ram[78]  = 1100001110110010;
    ram[79]  = 1010000111011001;
    ram[80]  = 1101000011101100;
    ram[81]  = 0101011110001001;
    ram[82]  = 1001010000111011;
    ram[83]  = 1100101000011101;
    ram[84]  = 1110010100001110;
    ram[85]  = 1011001010000111;
    ram[86]  = 0010011010111100;
    ram[87]  = 0001001101011110;
    ram[88]  = 1111011001010000;
    ram[89]  = 1011101100101000;
    ram[90]  = 0110001001101011;
    ram[91]  = 1000111011001010;
    ram[92]  = 1000011101100101;
    ram[93]  = 1100001110110010;
    ram[94]  = 0101111000100110;
    ram[95]  = 1101000011101100;
    ram[96]  = 1010100001110110;
    ram[97]  = 1001010000111011;
    ram[98]  = 0011010111100010;
    ram[99]  = 0001101011110001;
    ram[100] = 1011001010000111;
    ram[101] = 0010011010111100;
    ram[102] = 1110110010100001;
    ram[103] = 0000100110101111;
    ram[104] = 1011101100101000;
    ram[105] = 0110001001101011;
    ram[106] = 0111000100110101;
    ram[107] = 1000011101100101;
    ram[108] = 0011110001001101;
    ram[109] = 1010000111011001;
    ram[110] = 0010111100010011;
    ram[111] = 0101011110001001;
    ram[112] = 0110101111000100;
    ram[113] = 1100101000011101;
    ram[114] = 0001101011110001;
    ram[115] = 0100110101111000;
    ram[116] = 1101100101000011;
    ram[117] = 0001001101011110;
    ram[118] = 1111011001010000;
    ram[119] = 1011101100101000;
    ram[120] = 0110001001101011;
    ram[121] = 1000111011001010;
    ram[122] = 0111100010011010;
    ram[123] = 0011110001001101;
    ram[124] = 0101111000100110;
    ram[125] = 1101000011101100;
    ram[126] = 1010100001110110;
    ram[127] = 0110101111000100;
    ram[128] = 0011010111100010;
    ram[129] = 1110010100001110;
    ram[130] = 1011001010000111;
    ram[131] = 1101100101000011;
    ram[132] = 0001001101011110;
    ram[133] = 0000100110101111;
    ram[134] = 1011101100101000;
    ram[135] = 1001110110010100;
    ram[136] = 1000111011001010;
    ram[137] = 1000011101100101;
    ram[138] = 0011110001001101;
    ram[139] = 0101111000100110;
    ram[140] = 0010111100010011;
    ram[141] = 1010100001110110;
    ram[142] = 1001010000111011;
    ram[143] = 0011010111100010;
    ram[144] = 1110010100001110;
    ram[145] = 1011001010000111;
    ram[146] = 0010011010111100;
    ram[147] = 0001001101011110;
    ram[148] = 0000100110101111;
    ram[149] = 0100010011010111;
    ram[150] = 1001110110010100;
    ram[151] = 0111000100110101;
    ram[152] = 0111100010011010;
    ram[153] = 0011110001001101;
    ram[154] = 1010000111011001;
    ram[155] = 0010111100010011;
    ram[156] = 1010100001110110;
    ram[157] = 1001010000111011;
    ram[158] = 1100101000011101;
    ram[159] = 0001101011110001;
    ram[160] = 1011001010000111;
    ram[161] = 0010011010111100;
    ram[162] = 1110110010100001;
    ram[163] = 1111011001010000;
    ram[164] = 1011101100101000;
    ram[165] = 1001110110010100;
    ram[166] = 0111000100110101;
    ram[167] = 1000011101100101;
    ram[168] = 1100001110110010;
    ram[169] = 0101111000100110;
    ram[170] = 1101000011101100;
    ram[171] = 1010100001110110;
    ram[172] = 1001010000111011;
    ram[173] = 1100101000011101;
    ram[174] = 1110010100001110;
    ram[175] = 0100110101111000;
    ram[176] = 0010011010111100;
    ram[177] = 0001001101011110;
    ram[178] = 0000100110101111;
    ram[179] = 1011101100101000;
    ram[180] = 1001110110010100;
    ram[181] = 0111000100110101;
    ram[182] = 1000011101100101;
    ram[183] = 0011110001001101;
    ram[184] = 0101111000100110;
    ram[185] = 1101000011101100;
    ram[186] = 1010100001110110;
    ram[187] = 0110101111000100;
    ram[188] = 1100101000011101;
    ram[189] = 0001101011110001;
    ram[190] = 1011001010000111;
    ram[191] = 1101100101000011;
    ram[192] = 0001001101011110;
    ram[193] = 1111011001010000;
    ram[194] = 1011101100101000;
    ram[195] = 0110001001101011;
    ram[196] = 1000111011001010;
    ram[197] = 0111100010011010;
    ram[198] = 1100001110110010;
    ram[199] = 0101111000100110;
    ram[200] = 0010111100010011;
    ram[201] = 0101011110001001;
    ram[202] = 0110101111000100;
    ram[203] = 0011010111100010;
    ram[204] = 1110010100001110;
    ram[205] = 0100110101111000;
    ram[206] = 0010011010111100;
    ram[207] = 1110110010100001;
    ram[208] = 1111011001010000;
    ram[209] = 1011101100101000;
    ram[210] = 0110001001101011;
    ram[211] = 1000111011001010;
    ram[212] = 1000011101100101;
    ram[213] = 0011110001001101;
    ram[214] = 0101111000100110;
    ram[215] = 1101000011101100;
    ram[216] = 0101011110001001;
    ram[217] = 0110101111000100;
    ram[218] = 1100101000011101;
    ram[219] = 0001101011110001;
    ram[220] = 0100110101111000;
    ram[221] = 1101100101000011;
    ram[222] = 1110110010100001;
    ram[223] = 0000100110101111;
    ram[224] = 0100010011010111;
    ram[225] = 0110001001101011;
    ram[226] = 0111000100110101;
    ram[227] = 0111100010011010;
    ram[228] = 0011110001001101;
    ram[229] = 1010000111011001;
    ram[230] = 1101000011101100;
    ram[231] = 1010100001110110;
    ram[232] = 0110101111000100;
    ram[233] = 1100101000011101;
    ram[234] = 0001101011110001;
    ram[235] = 0100110101111000;
    ram[236] = 1101100101000011;
    ram[237] = 0001001101011110;
    ram[238] = 0000100110101111;
    ram[239] = 0100010011010111;
    ram[240] = 1001110110010100;
    ram[241] = 1000111011001010;
    ram[242] = 1000011101100101;
    ram[243] = 0011110001001101;
    ram[244] = 0101111000100110;
    ram[245] = 0010111100010011;
    ram[246] = 1010100001110110;
    ram[247] = 0110101111000100;
    ram[248] = 0011010111100010;
    ram[249] = 0001101011110001;
    ram[250] = 0100110101111000;
    ram[251] = 0010011010111100;
    ram[252] = 0001001101011110;
    ram[253] = 0000100110101111;
    ram[254] = 1011101100101000;
  end
  
  always @(posedge clk) begin 
   if (ena) begin
      if (wea)
          ram[addra] <= dia;
   end
  end
    
  always @(posedge clk) begin 
    if (enb)
      dob <= ram[addrb];
  end
  
endmodule

//MODULE OBTAINED ON THE XILINX WEBSITE